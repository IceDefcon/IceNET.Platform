library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity temp is
port
(    
    clock : in std_logic;
    reset : in std_logic;

    input : in std_logic;
    output : out std_logic
);
end temp;

architecture rtl of temp is

--
-- CODE
--

end rtl;